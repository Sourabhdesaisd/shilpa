module ex_mem_pipeline (
    input  wire        clk,
    input  wire        rst,

    // Inputs from EX stage
    input  wire [31:0] ex_result_in,
    input  wire [31:0] addr_result_in,
    input  wire [4:0]  rd_in,
    input  wire        mwr_in,
    input  wire        werf_in,
    input  wire        b_mux_in,
    input  wire wb_sel_in,
    

    // Outputs to MEM stage
    output reg  [31:0] ex_result_out,
    output reg  [31:0] addr_result_out,
    output reg  [4:0]  rd_out,
    output reg         mwr_out,
    output reg         werf_out,
    output reg         b_mux_out,
    output reg  wb_sel_out
    
);

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            ex_result_out   <= 32'b0;
            addr_result_out <= 32'b0;
            rd_out          <= 5'b0;
            mwr_out         <= 1'b0;
            werf_out        <= 1'b0;
            b_mux_out       <= 1'b0;
            wb_sel_out <= 1'b0;
            
        end 
        else begin
            ex_result_out   <= ex_result_in;
            addr_result_out <= addr_result_in;
            rd_out          <= rd_in;
            mwr_out         <= mwr_in;
            werf_out        <= werf_in;
            b_mux_out       <= b_mux_in;
            wb_sel_out <= wb_sel_in;
            
        end
    end

endmodule
